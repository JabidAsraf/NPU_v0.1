`timescale 1ns/1ps // time_unit/time_precision

`define FP32

`ifdef FP32
    `define MODE 1
    `define MULTIPLIER_UNIT fp32_multiplier
    `define NURON_WIDTH 32
    `define CONV_F2B_FUNC $shortrealtobits
    `define CONV_B2F_FUNC $bitstoshortreal
`else
    `define MODE 0
    `define MULTIPLIER_UNIT fp16_multiplier
    `define NURON_WIDTH 16
    `define CONV_F2B_FUNC float2bin
    `define CONV_B2F_FUNC bin2float
`endif

module tb_fm_err_chk_ind;
  
    reg                     clk;
    reg                     reset_b;
    reg  [`NURON_WIDTH-1:0] a;
    reg  [`NURON_WIDTH-1:0] b;
    reg                     start;
    reg                     clear;
    wire                    valid;
    wire [`NURON_WIDTH-1:0] out; 
      
    shortreal i, j;
    shortreal max_err = 0;
    shortreal min_err = 0;

    int f_handle;
    int info_f_handle;
    int count;

    `MULTIPLIER_UNIT dut
    (
        .clk     ( clk     ),
        .reset_b ( reset_b ),
        .input_a ( a       ),
        .input_b ( b       ),
        .start   ( start   ),
        .clear   ( clear   ),
        .valid   ( valid   ),
        .result  ( out     )
    );


    initial begin
        clk <= 0;
        forever #0.5 clk <= ~clk;
    end
    

    initial begin
        $write("%c[1;34m",27);
   
        $display("Runnning multiplier error check test in %0s mode", (`MODE ? "FP32" : "FP16") );

        reset();

        multi_op(99.99, 13);
        
        $write("%c[0m",27);
    
        #20 $stop;
    end
    

    task reset();
        reset_b   <=  1'b0;
        a         <=  `NURON_WIDTH'd0;
        b         <=  `NURON_WIDTH'd0;
        start     <=  1'b0;
        clear     <=  1'b0;
        count     <=  0;
        @(posedge clk) reset_b <= 1'b1;
    endtask
    

    task multi_op(shortreal float_a, shortreal float_b);
        shortreal exp, act, err, err_per;

        exp        = 0;
        act        = 0;
        err        = 0;
        err_per    = 0;

        a         <=  `CONV_F2B_FUNC(float_a);
        b         <=  `CONV_F2B_FUNC(float_b);
        @(posedge clk) start <= 1'b1;
        @(posedge clk) start <= 1'b0;
        wait(valid);
        @(posedge clk) clear <= 1'b1;
        @(posedge clk) clear <= 1'b0;
        
        exp     = (float_a*float_b);
        act     = `CONV_B2F_FUNC(out);
        err     = (exp > act) ? (exp - act) : (act - exp);

        if(((float_a*float_b) > 0.0001) || ((float_a*float_b) < -0.0001)) begin
            err_per = (exp == 0)  ? 0 : (err/exp)*100;
        end else begin
            err_per = 0;
        end

        if(max_err < err_per) begin
            max_err = err_per;
        end

        if(min_err > err_per) begin
            min_err = err_per;
        end

        `ifndef FP32
        
            count = count + 1;
            $display("[%20t] :: Multiplication number: %0d", $time, count);
            
            $display("-------------------------------------------------------------------------------------------------------------");
            $display("input a in binary         = %16b :: input a in float         = %0f",   a,              float_a );
            $display("input b in binary         = %16b :: input b in float         = %0f",   b,              float_b );
            
            $display("mantisa[10:0]             = %11b                                  ",   dut.mantisa             );
            $display("mantisa_temp[10:0]        = %11b                                  ",   dut.mantisa_temp        );
            $display("exponent[4:0]             = %5b                                   ",   dut.exponent            );
            $display("ovcheck                   = %1b                                   ",   dut.ovcheck             );
            $display("elcheck                   = %1b                                   ",   dut.elcheck             );
            $display("zcheck                    = %1b                                   ",   dut.zcheck              );
            $display("mantisa_pre_el[9:0]       = %10b                                  ",   dut.mantisa_pre_el      );
            $display("mantisa_final[9:0]        = %10b                                  ",   dut.mantisa_final       );
            $display("exponent_final[4:0]       = %5b                                   ",   dut.exponent_final      );
            
            $display("expected output in binary = %16b :: expected output in float = %0f",   float2bin(exp), exp     );
            $display("actual output in binary   = %16b :: actual output in float   = %0f\n", out,            act     );
            $display("error absolute            = %0f",                                      err                     );    
            $display("error percentage          = %0f",                                      err_per                 );    
            $display("-------------------------------------------------------------------------------------------------------------\n\n");
        
        `else
            
            count = count + 1;
            $display("[%20t] :: Multiplication number: %0d", $time, count);
            
            $display("-------------------------------------------------------------------------------------------------------------");
            $display("input a in binary         = %32b :: input a in float         = %0f",   a,                     float_a );
            $display("input b in binary         = %32b :: input b in float         = %0f",   b,                     float_b );
                        
            $display("expected output in binary = %32b :: expected output in float = %0f",   $shortrealtobits(exp), exp     );
            $display("actual output in binary   = %32b :: actual output in float   = %0f\n", out,                   act     );
            $display("error absolute            = %0f",                                      err                            );    
            $display("error percentage          = %0f",                                      err_per                        );    
            $display("-------------------------------------------------------------------------------------------------------------\n\n");
        
        `endif
    endtask
      

    function [15:0] float2bin (shortreal float_a);
        logic [31:0] fp32;
        logic [7:0]  exp_temp;
        logic [22:0] man_temp;
        fp32     [31:0] = $shortrealtobits(float_a);
        exp_temp [7:0]  = ((fp32[30:23] - 8'd127) <= (-15)) && (float_a < 1) && (float_a > -1) ? 0                    : (fp32[30:23] - 8'd127 + 8'd15);
        man_temp [22:0] = ((fp32[30:23] - 8'd127) == (-15))                  ? {1'b1,fp32[22:1]}    : 
                          ((fp32[30:23] - 8'd127) == (-16))                  ? {2'b01, fp32[22:2]}  : 
                          ((fp32[30:23] - 8'd127) == (-17))                  ? {3'b001, fp32[22:3]} : fp32[22:0];
        return ((float_a == 0) ? 16'd0 : {fp32[31], exp_temp[4:0], man_temp[22:13]});
    endfunction
    

    function shortreal bin2float (logic [15:0] fp16);
        logic [31:0] fp32;
        logic [7:0]  exp_temp;
        logic [22:0] man_temp;
    
        exp_temp [7:0]  = {3'd0, fp16[14:10]} - 8'd15 + 8'd127;
        man_temp [22:0] = {fp16[9:0],13'd0};
        fp32     [31:0] = {fp16[15], exp_temp[7:0], man_temp[22:0]};
    
        return (~(|fp16[15:0]) ? 0 : $bitstoshortreal(fp32[31:0]));
    endfunction
  

endmodule
